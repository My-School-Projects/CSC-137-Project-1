// atter_test.v

module adder_test(cin, a, b, s, cout);

    output reg cin;
    output reg [3:0] a, b;

    input [3:0] s;
    input cout;

    initial begin

        $monitor("a %b cin  %b\nb %b cout %b\ns %b\n", a, cin, b, cout, s);

        cin = 0;
        a = 4'b0000;
        b = 4'b0000;

        #10

        a = 4'b0000;
        b = 4'b0001;

        #10

        a = 4'b0000;
        b = 4'b0010;

        #10

        a = 4'b0000;
        b = 4'b0011;

        #10

        a = 4'b0000;
        b = 4'b0100;

        #10

        a = 4'b0000;
        b = 4'b0101;

        #10

        a = 4'b0000;
        b = 4'b0110;

        #10

        a = 4'b0000;
        b = 4'b0111;

        #10

        a = 4'b0000;
        b = 4'b1000;

        #10

        a = 4'b0000;
        b = 4'b1001;

        #10

        a = 4'b0000;
        b = 4'b1010;

        #10

        a = 4'b0000;
        b = 4'b1011;

        #10

        a = 4'b0000;
        b = 4'b1100;

        #10

        a = 4'b0000;
        b = 4'b1101;

        #10

        a = 4'b0000;
        b = 4'b1110;

        #10

        a = 4'b0000;
        b = 4'b1111;

        #10

        a = 4'b0001;
        b = 4'b0000;

        #10

        a = 4'b0001;
        b = 4'b0001;

        #10

        a = 4'b0001;
        b = 4'b0010;

        #10

        a = 4'b0001;
        b = 4'b0011;

        #10

        a = 4'b0001;
        b = 4'b0100;

        #10

        a = 4'b0001;
        b = 4'b0101;

        #10

        a = 4'b0001;
        b = 4'b0110;

        #10

        a = 4'b0001;
        b = 4'b0111;

        #10

        a = 4'b0001;
        b = 4'b1000;

        #10

        a = 4'b0001;
        b = 4'b1001;

        #10

        a = 4'b0001;
        b = 4'b1010;

        #10

        a = 4'b0001;
        b = 4'b1011;

        #10

        a = 4'b0001;
        b = 4'b1100;

        #10

        a = 4'b0001;
        b = 4'b1101;

        #10

        a = 4'b0001;
        b = 4'b1110;

        #10

        a = 4'b0001;
        b = 4'b1111;

        #10

        a = 4'b0010;
        b = 4'b0000;

        #10

        a = 4'b0010;
        b = 4'b0001;

        #10

        a = 4'b0010;
        b = 4'b0010;

        #10

        a = 4'b0010;
        b = 4'b0011;

        #10

        a = 4'b0010;
        b = 4'b0100;

        #10

        a = 4'b0010;
        b = 4'b0101;

        #10

        a = 4'b0010;
        b = 4'b0110;

        #10

        a = 4'b0010;
        b = 4'b0111;

        #10

        a = 4'b0010;
        b = 4'b1000;

        #10

        a = 4'b0010;
        b = 4'b1001;

        #10

        a = 4'b0010;
        b = 4'b1010;

        #10

        a = 4'b0010;
        b = 4'b1011;

        #10

        a = 4'b0010;
        b = 4'b1100;

        #10

        a = 4'b0010;
        b = 4'b1101;

        #10

        a = 4'b0010;
        b = 4'b1110;

        #10

        a = 4'b0010;
        b = 4'b1111;

        #10

        a = 4'b0011;
        b = 4'b0000;

        #10

        a = 4'b0011;
        b = 4'b0001;

        #10

        a = 4'b0011;
        b = 4'b0010;

        #10

        a = 4'b0011;
        b = 4'b0011;

        #10

        a = 4'b0011;
        b = 4'b0100;

        #10

        a = 4'b0011;
        b = 4'b0101;

        #10

        a = 4'b0011;
        b = 4'b0110;

        #10

        a = 4'b0011;
        b = 4'b0111;

        #10

        a = 4'b0011;
        b = 4'b1000;

        #10

        a = 4'b0011;
        b = 4'b1001;

        #10

        a = 4'b0011;
        b = 4'b1010;

        #10

        a = 4'b0011;
        b = 4'b1011;

        #10

        a = 4'b0011;
        b = 4'b1100;

        #10

        a = 4'b0011;
        b = 4'b1101;

        #10

        a = 4'b0011;
        b = 4'b1110;

        #10

        a = 4'b0011;
        b = 4'b1111;

        #10

        a = 4'b0100;
        b = 4'b0000;

        #10

        a = 4'b0100;
        b = 4'b0001;

        #10

        a = 4'b0100;
        b = 4'b0010;

        #10

        a = 4'b0100;
        b = 4'b0011;

        #10

        a = 4'b0100;
        b = 4'b0100;

        #10

        a = 4'b0100;
        b = 4'b0101;

        #10

        a = 4'b0100;
        b = 4'b0110;

        #10

        a = 4'b0100;
        b = 4'b0111;

        #10

        a = 4'b0100;
        b = 4'b1000;

        #10

        a = 4'b0100;
        b = 4'b1001;

        #10

        a = 4'b0100;
        b = 4'b1010;

        #10

        a = 4'b0100;
        b = 4'b1011;

        #10

        a = 4'b0100;
        b = 4'b1100;

        #10

        a = 4'b0100;
        b = 4'b1101;

        #10

        a = 4'b0100;
        b = 4'b1110;

        #10

        a = 4'b0100;
        b = 4'b1111;

        #10

        a = 4'b0101;
        b = 4'b0000;

        #10

        a = 4'b0101;
        b = 4'b0001;

        #10

        a = 4'b0101;
        b = 4'b0010;

        #10

        a = 4'b0101;
        b = 4'b0011;

        #10

        a = 4'b0101;
        b = 4'b0100;

        #10

        a = 4'b0101;
        b = 4'b0101;

        #10

        a = 4'b0101;
        b = 4'b0110;

        #10

        a = 4'b0101;
        b = 4'b0111;

        #10

        a = 4'b0101;
        b = 4'b1000;

        #10

        a = 4'b0101;
        b = 4'b1001;

        #10

        a = 4'b0101;
        b = 4'b1010;

        #10

        a = 4'b0101;
        b = 4'b1011;

        #10

        a = 4'b0101;
        b = 4'b1100;

        #10

        a = 4'b0101;
        b = 4'b1101;

        #10

        a = 4'b0101;
        b = 4'b1110;

        #10

        a = 4'b0101;
        b = 4'b1111;

        #10

        a = 4'b0110;
        b = 4'b0000;

        #10

        a = 4'b0110;
        b = 4'b0001;

        #10

        a = 4'b0110;
        b = 4'b0010;

        #10

        a = 4'b0110;
        b = 4'b0011;

        #10

        a = 4'b0110;
        b = 4'b0100;

        #10

        a = 4'b0110;
        b = 4'b0101;

        #10

        a = 4'b0110;
        b = 4'b0110;

        #10

        a = 4'b0110;
        b = 4'b0111;

        #10

        a = 4'b0110;
        b = 4'b1000;

        #10

        a = 4'b0110;
        b = 4'b1001;

        #10

        a = 4'b0110;
        b = 4'b1010;

        #10

        a = 4'b0110;
        b = 4'b1011;

        #10

        a = 4'b0110;
        b = 4'b1100;

        #10

        a = 4'b0110;
        b = 4'b1101;

        #10

        a = 4'b0110;
        b = 4'b1110;

        #10

        a = 4'b0110;
        b = 4'b1111;

        #10

        a = 4'b0111;
        b = 4'b0000;

        #10

        a = 4'b0111;
        b = 4'b0001;

        #10

        a = 4'b0111;
        b = 4'b0010;

        #10

        a = 4'b0111;
        b = 4'b0011;

        #10

        a = 4'b0111;
        b = 4'b0100;

        #10

        a = 4'b0111;
        b = 4'b0101;

        #10

        a = 4'b0111;
        b = 4'b0110;

        #10

        a = 4'b0111;
        b = 4'b0111;

        #10

        a = 4'b0111;
        b = 4'b1000;

        #10

        a = 4'b0111;
        b = 4'b1001;

        #10

        a = 4'b0111;
        b = 4'b1010;

        #10

        a = 4'b0111;
        b = 4'b1011;

        #10

        a = 4'b0111;
        b = 4'b1100;

        #10

        a = 4'b0111;
        b = 4'b1101;

        #10

        a = 4'b0111;
        b = 4'b1110;

        #10

        a = 4'b0111;
        b = 4'b1111;

        #10

        a = 4'b1000;
        b = 4'b0000;

        #10

        a = 4'b1000;
        b = 4'b0001;

        #10

        a = 4'b1000;
        b = 4'b0010;

        #10

        a = 4'b1000;
        b = 4'b0011;

        #10

        a = 4'b1000;
        b = 4'b0100;

        #10

        a = 4'b1000;
        b = 4'b0101;

        #10

        a = 4'b1000;
        b = 4'b0110;

        #10

        a = 4'b1000;
        b = 4'b0111;

        #10

        a = 4'b1000;
        b = 4'b1000;

        #10

        a = 4'b1000;
        b = 4'b1001;

        #10

        a = 4'b1000;
        b = 4'b1010;

        #10

        a = 4'b1000;
        b = 4'b1011;

        #10

        a = 4'b1000;
        b = 4'b1100;

        #10

        a = 4'b1000;
        b = 4'b1101;

        #10

        a = 4'b1000;
        b = 4'b1110;

        #10

        a = 4'b1000;
        b = 4'b1111;

        #10

        a = 4'b1001;
        b = 4'b0000;

        #10

        a = 4'b1001;
        b = 4'b0001;

        #10

        a = 4'b1001;
        b = 4'b0010;

        #10

        a = 4'b1001;
        b = 4'b0011;

        #10

        a = 4'b1001;
        b = 4'b0100;

        #10

        a = 4'b1001;
        b = 4'b0101;

        #10

        a = 4'b1001;
        b = 4'b0110;

        #10

        a = 4'b1001;
        b = 4'b0111;

        #10

        a = 4'b1001;
        b = 4'b1000;

        #10

        a = 4'b1001;
        b = 4'b1001;

        #10

        a = 4'b1001;
        b = 4'b1010;

        #10

        a = 4'b1001;
        b = 4'b1011;

        #10

        a = 4'b1001;
        b = 4'b1100;

        #10

        a = 4'b1001;
        b = 4'b1101;

        #10

        a = 4'b1001;
        b = 4'b1110;

        #10

        a = 4'b1001;
        b = 4'b1111;

        #10

        a = 4'b1010;
        b = 4'b0000;

        #10

        a = 4'b1010;
        b = 4'b0001;

        #10

        a = 4'b1010;
        b = 4'b0010;

        #10

        a = 4'b1010;
        b = 4'b0011;

        #10

        a = 4'b1010;
        b = 4'b0100;

        #10

        a = 4'b1010;
        b = 4'b0101;

        #10

        a = 4'b1010;
        b = 4'b0110;

        #10

        a = 4'b1010;
        b = 4'b0111;

        #10

        a = 4'b1010;
        b = 4'b1000;

        #10

        a = 4'b1010;
        b = 4'b1001;

        #10

        a = 4'b1010;
        b = 4'b1010;

        #10

        a = 4'b1010;
        b = 4'b1011;

        #10

        a = 4'b1010;
        b = 4'b1100;

        #10

        a = 4'b1010;
        b = 4'b1101;

        #10

        a = 4'b1010;
        b = 4'b1110;

        #10

        a = 4'b1010;
        b = 4'b1111;

        #10

        a = 4'b1011;
        b = 4'b0000;

        #10

        a = 4'b1011;
        b = 4'b0001;

        #10

        a = 4'b1011;
        b = 4'b0010;

        #10

        a = 4'b1011;
        b = 4'b0011;

        #10

        a = 4'b1011;
        b = 4'b0100;

        #10

        a = 4'b1011;
        b = 4'b0101;

        #10

        a = 4'b1011;
        b = 4'b0110;

        #10

        a = 4'b1011;
        b = 4'b0111;

        #10

        a = 4'b1011;
        b = 4'b1000;

        #10

        a = 4'b1011;
        b = 4'b1001;

        #10

        a = 4'b1011;
        b = 4'b1010;

        #10

        a = 4'b1011;
        b = 4'b1011;

        #10

        a = 4'b1011;
        b = 4'b1100;

        #10

        a = 4'b1011;
        b = 4'b1101;

        #10

        a = 4'b1011;
        b = 4'b1110;

        #10

        a = 4'b1011;
        b = 4'b1111;

        #10

        a = 4'b1100;
        b = 4'b0000;

        #10

        a = 4'b1100;
        b = 4'b0001;

        #10

        a = 4'b1100;
        b = 4'b0010;

        #10

        a = 4'b1100;
        b = 4'b0011;

        #10

        a = 4'b1100;
        b = 4'b0100;

        #10

        a = 4'b1100;
        b = 4'b0101;

        #10

        a = 4'b1100;
        b = 4'b0110;

        #10

        a = 4'b1100;
        b = 4'b0111;

        #10

        a = 4'b1100;
        b = 4'b1000;

        #10

        a = 4'b1100;
        b = 4'b1001;

        #10

        a = 4'b1100;
        b = 4'b1010;

        #10

        a = 4'b1100;
        b = 4'b1011;

        #10

        a = 4'b1100;
        b = 4'b1100;

        #10

        a = 4'b1100;
        b = 4'b1101;

        #10

        a = 4'b1100;
        b = 4'b1110;

        #10

        a = 4'b1100;
        b = 4'b1111;

        #10

        a = 4'b1101;
        b = 4'b0000;

        #10

        a = 4'b1101;
        b = 4'b0001;

        #10

        a = 4'b1101;
        b = 4'b0010;

        #10

        a = 4'b1101;
        b = 4'b0011;

        #10

        a = 4'b1101;
        b = 4'b0100;

        #10

        a = 4'b1101;
        b = 4'b0101;

        #10

        a = 4'b1101;
        b = 4'b0110;

        #10

        a = 4'b1101;
        b = 4'b0111;

        #10

        a = 4'b1101;
        b = 4'b1000;

        #10

        a = 4'b1101;
        b = 4'b1001;

        #10

        a = 4'b1101;
        b = 4'b1010;

        #10

        a = 4'b1101;
        b = 4'b1011;

        #10

        a = 4'b1101;
        b = 4'b1100;

        #10

        a = 4'b1101;
        b = 4'b1101;

        #10

        a = 4'b1101;
        b = 4'b1110;

        #10

        a = 4'b1101;
        b = 4'b1111;

        #10

        a = 4'b1110;
        b = 4'b0000;

        #10

        a = 4'b1110;
        b = 4'b0001;

        #10

        a = 4'b1110;
        b = 4'b0010;

        #10

        a = 4'b1110;
        b = 4'b0011;

        #10

        a = 4'b1110;
        b = 4'b0100;

        #10

        a = 4'b1110;
        b = 4'b0101;

        #10

        a = 4'b1110;
        b = 4'b0110;

        #10

        a = 4'b1110;
        b = 4'b0111;

        #10

        a = 4'b1110;
        b = 4'b1000;

        #10

        a = 4'b1110;
        b = 4'b1001;

        #10

        a = 4'b1110;
        b = 4'b1010;

        #10

        a = 4'b1110;
        b = 4'b1011;

        #10

        a = 4'b1110;
        b = 4'b1100;

        #10

        a = 4'b1110;
        b = 4'b1101;

        #10

        a = 4'b1110;
        b = 4'b1110;

        #10

        a = 4'b1110;
        b = 4'b1111;

        #10

        a = 4'b1111;
        b = 4'b0000;

        #10

        a = 4'b1111;
        b = 4'b0001;

        #10

        a = 4'b1111;
        b = 4'b0010;

        #10

        a = 4'b1111;
        b = 4'b0011;

        #10

        a = 4'b1111;
        b = 4'b0100;

        #10

        a = 4'b1111;
        b = 4'b0101;

        #10

        a = 4'b1111;
        b = 4'b0110;

        #10

        a = 4'b1111;
        b = 4'b0111;

        #10

        a = 4'b1111;
        b = 4'b1000;

        #10

        a = 4'b1111;
        b = 4'b1001;

        #10

        a = 4'b1111;
        b = 4'b1010;

        #10

        a = 4'b1111;
        b = 4'b1011;

        #10

        a = 4'b1111;
        b = 4'b1100;

        #10

        a = 4'b1111;
        b = 4'b1101;

        #10

        a = 4'b1111;
        b = 4'b1110;

        #10

        a = 4'b1111;
        b = 4'b1111;

        $finish;

    end

endmodule

module adder_bench();

    wire cin, cout;
    wire [3:0] a, b, s;

    adder u(cin, a, b, s, cout);

    adder_test t(cin, a, b, s, cout);

endmodule
