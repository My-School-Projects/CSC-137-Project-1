module pgu (
    a0,
    a1,
    a2,
    a3,
    b0,
    b1,
    b2,
    b3,
    p0,
    p1,
    p2,
    p3,
    g0,
    g1,
    g2,
    g3
)

input a0;
input a1;
input a2;
input a3;
input b0;
input b1;
input b2;
input b3;

output p0;
output p1;
output p2;
output p3;
output g0;
output g1;
output g2;
output g3;